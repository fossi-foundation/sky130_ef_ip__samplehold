magic
tech sky130A
magscale 1 2
timestamp 1750254930
<< dnwell >>
rect 373 -3022 2461 2010
<< nwell >>
rect 264 1804 2570 2130
rect 264 782 579 1804
rect 2255 782 2570 1804
rect 264 673 2570 782
rect 264 -1800 614 673
rect 1957 -297 2570 673
rect 2240 -1800 2570 -297
rect 264 -2816 579 -1800
rect 2255 -2816 2570 -1800
rect 264 -3133 2570 -2816
<< mvpsubdiff >>
rect 1786 874 1806 1236
<< mvnsubdiff >>
rect 330 2044 2504 2064
rect 330 2010 410 2044
rect 2424 2010 2504 2044
rect 330 1990 2504 2010
rect 330 1984 404 1990
rect 330 -2985 350 1984
rect 384 -2985 404 1984
rect 2430 1984 2504 1990
rect 330 -2991 404 -2985
rect 2430 -2985 2450 1984
rect 2484 -2985 2504 1984
rect 2430 -2991 2504 -2985
rect 330 -3011 2504 -2991
rect 330 -3045 410 -3011
rect 2424 -3045 2504 -3011
rect 330 -3065 2504 -3045
<< mvnsubdiffcont >>
rect 410 2010 2424 2044
rect 350 -2985 384 1984
rect 2450 -2985 2484 1984
rect 410 -3045 2424 -3011
<< locali >>
rect 350 2010 410 2044
rect 2424 2010 2484 2044
rect 350 1984 2484 2010
rect 384 1921 2450 1984
rect 384 782 534 1921
rect 579 856 768 1676
rect 1169 1655 1343 1677
rect 1169 974 1221 1655
rect 1297 974 1343 1655
rect 1169 856 1343 974
rect 1753 1657 2282 1677
rect 1753 976 1802 1657
rect 1878 1147 2282 1657
rect 1878 1146 1927 1147
rect 1878 976 1882 1146
rect 1753 856 1882 976
rect 2130 856 2282 1147
rect 2352 782 2450 1921
rect 384 642 2450 782
rect 384 -158 712 642
rect 1870 -158 2450 642
rect 384 -185 2450 -158
rect 384 -358 500 -185
rect 2364 -358 2450 -185
rect 384 -374 2450 -358
rect 384 -1694 712 -374
rect 2140 -1694 2450 -374
rect 384 -1788 2450 -1694
rect 384 -2628 491 -1788
rect 562 -1955 2262 -1866
rect 562 -2670 714 -1955
rect 2120 -2670 2262 -1955
rect 2329 -2621 2450 -1788
rect 434 -2711 2405 -2670
rect 434 -2881 545 -2711
rect 2354 -2881 2405 -2711
rect 434 -2943 2405 -2881
rect 350 -3011 384 -2985
rect 2450 -3011 2484 -2985
rect 350 -3045 410 -3011
rect 2424 -3045 2484 -3011
<< viali >>
rect 1221 974 1297 1655
rect 1802 976 1878 1657
rect 500 -358 2364 -185
rect 545 -2881 2354 -2711
<< metal1 >>
rect 393 1841 2463 1863
rect 393 1622 544 1841
rect 842 1657 2463 1841
rect 842 1655 1802 1657
rect 842 1622 1221 1655
rect 393 1606 1221 1622
rect 824 1098 888 1606
rect 340 919 540 990
rect 943 919 980 1531
rect 340 867 894 919
rect 972 867 980 919
rect 340 790 540 867
rect 943 701 980 867
rect 1052 802 1101 1472
rect 1211 974 1221 1606
rect 1297 1606 1802 1655
rect 1297 974 1308 1606
rect 1406 1096 1470 1606
rect 1211 959 1308 974
rect 1534 802 1571 1532
rect 1052 753 1571 802
rect 909 664 1099 701
rect 909 500 946 664
rect 1062 500 1099 664
rect 793 438 866 453
rect 793 -46 803 438
rect 857 -46 866 438
rect 793 -59 866 -46
rect 964 -92 1036 456
rect 1158 439 1207 753
rect 1534 701 1571 753
rect 1620 800 1669 1471
rect 1791 976 1802 1606
rect 1878 1606 2463 1657
rect 1878 976 1888 1606
rect 1791 964 1888 976
rect 1961 919 2032 1039
rect 1961 861 2032 867
rect 1620 751 1792 800
rect 1490 664 1680 701
rect 1490 500 1527 664
rect 1643 500 1680 664
rect 1201 -45 1207 439
rect 1158 -57 1207 -45
rect 1375 440 1448 451
rect 1375 -44 1382 440
rect 1436 -44 1448 440
rect 1375 -61 1448 -44
rect 1552 -92 1624 451
rect 1743 440 1792 751
rect 1786 -44 1792 440
rect 1743 -59 1792 -44
rect 326 -185 2478 -92
rect 326 -358 500 -185
rect 2364 -358 2478 -185
rect 326 -368 2478 -358
rect 904 -449 959 -397
rect 1040 -449 1046 -397
rect 904 -453 1046 -449
rect 745 -1042 867 -1036
rect 745 -1197 751 -1042
rect 333 -1395 751 -1197
rect 860 -1395 867 -1042
rect 333 -1397 867 -1395
rect 745 -1405 867 -1397
rect 904 -1667 939 -453
rect 1370 -455 1376 -402
rect 1457 -455 1525 -402
rect 1370 -458 1525 -455
rect 1190 -501 1292 -495
rect 1190 -885 1196 -501
rect 1286 -885 1292 -501
rect 1190 -891 1292 -885
rect 977 -1041 1099 -1035
rect 977 -1394 984 -1041
rect 1093 -1394 1099 -1041
rect 977 -1400 1099 -1394
rect 1350 -1414 1356 -1048
rect 1446 -1414 1452 -1048
rect 1489 -1549 1525 -458
rect 1562 -501 1664 -495
rect 1562 -885 1568 -501
rect 1658 -885 1664 -501
rect 1755 -511 1876 -505
rect 1755 -864 1761 -511
rect 1870 -864 1876 -511
rect 1755 -870 1876 -864
rect 1988 -511 2109 -505
rect 1988 -864 1994 -511
rect 2103 -864 2109 -511
rect 1988 -870 2109 -864
rect 1562 -891 1664 -885
rect 2209 -1396 2526 -1196
rect 2209 -1402 2393 -1396
rect 1334 -1579 1685 -1549
rect 1334 -1585 1623 -1579
rect 1617 -1639 1623 -1585
rect 1679 -1639 1685 -1579
rect 1913 -1667 1948 -1460
rect 904 -1715 1948 -1667
rect 1051 -1845 1128 -1837
rect 1051 -1907 1128 -1901
rect 1051 -2031 1087 -1907
rect 887 -2067 1087 -2031
rect 1479 -2034 1515 -1715
rect 1728 -1845 1805 -1839
rect 1728 -1909 1805 -1901
rect 740 -2118 856 -2112
rect 740 -2255 746 -2118
rect 850 -2255 856 -2118
rect 740 -2261 856 -2255
rect 887 -2584 923 -2067
rect 1322 -2070 1515 -2034
rect 1756 -2032 1792 -1909
rect 2209 -2026 2217 -1402
rect 2387 -2026 2393 -1402
rect 1756 -2068 1949 -2032
rect 2209 -2036 2393 -2026
rect 967 -2118 1083 -2112
rect 967 -2255 973 -2118
rect 1077 -2255 1083 -2118
rect 967 -2261 1083 -2255
rect 1323 -2128 1440 -2122
rect 1323 -2252 1329 -2128
rect 1434 -2252 1440 -2128
rect 1323 -2258 1440 -2252
rect 1166 -2357 1282 -2351
rect 1166 -2494 1172 -2357
rect 1276 -2494 1282 -2357
rect 1166 -2500 1282 -2494
rect 1479 -2543 1515 -2070
rect 1552 -2357 1668 -2351
rect 1552 -2494 1558 -2357
rect 1662 -2494 1668 -2357
rect 1552 -2500 1668 -2494
rect 1750 -2357 1866 -2351
rect 1750 -2494 1756 -2357
rect 1860 -2494 1866 -2357
rect 1750 -2500 1866 -2494
rect 1347 -2579 1515 -2543
rect 1910 -2586 1946 -2068
rect 1978 -2357 2094 -2351
rect 1978 -2494 1984 -2357
rect 2088 -2494 2094 -2357
rect 1978 -2500 2094 -2494
rect 328 -2679 2515 -2670
rect 328 -2898 542 -2679
rect 840 -2711 2515 -2679
rect 2354 -2881 2515 -2711
rect 840 -2898 2515 -2881
rect 328 -2905 2515 -2898
<< via1 >>
rect 544 1622 842 1841
rect 894 867 972 919
rect 803 -46 857 438
rect 1961 867 2032 919
rect 1147 -45 1201 439
rect 1382 -44 1436 440
rect 1732 -44 1786 440
rect 959 -449 1040 -397
rect 751 -1395 860 -1042
rect 1376 -455 1457 -402
rect 1196 -885 1286 -501
rect 984 -1394 1093 -1041
rect 1356 -1414 1446 -1048
rect 1568 -885 1658 -501
rect 1761 -864 1870 -511
rect 1994 -864 2103 -511
rect 1623 -1639 1679 -1579
rect 1051 -1901 1128 -1845
rect 1728 -1901 1805 -1845
rect 746 -2255 850 -2118
rect 2217 -2026 2387 -1402
rect 973 -2255 1077 -2118
rect 1329 -2252 1434 -2128
rect 1172 -2494 1276 -2357
rect 1558 -2494 1662 -2357
rect 1756 -2494 1860 -2357
rect 1984 -2494 2088 -2357
rect 542 -2711 840 -2679
rect 542 -2881 545 -2711
rect 545 -2881 840 -2711
rect 542 -2898 840 -2881
<< metal2 >>
rect 529 1841 867 1856
rect 529 1622 544 1841
rect 842 1622 867 1841
rect 529 1606 867 1622
rect 529 -2670 660 1606
rect 886 867 894 919
rect 972 867 1961 919
rect 2032 867 2039 919
rect 795 439 1207 441
rect 795 438 1147 439
rect 795 -46 803 438
rect 857 -45 1147 438
rect 1201 -45 1207 439
rect 857 -46 1207 -45
rect 795 -47 1207 -46
rect 1376 440 1792 442
rect 1376 -44 1382 440
rect 1436 -44 1732 440
rect 1786 -44 1792 440
rect 1376 -46 1792 -44
rect 959 -397 1040 -47
rect 959 -455 1040 -449
rect 1376 -402 1457 -46
rect 1376 -461 1457 -455
rect 736 -501 2393 -489
rect 736 -885 1196 -501
rect 1286 -885 1568 -501
rect 1658 -511 2393 -501
rect 1658 -864 1761 -511
rect 1870 -864 1994 -511
rect 2103 -864 2393 -511
rect 1658 -885 2393 -864
rect 736 -893 2393 -885
rect 732 -1041 2127 -1034
rect 732 -1042 984 -1041
rect 732 -1395 751 -1042
rect 860 -1394 984 -1042
rect 1093 -1048 2127 -1041
rect 1093 -1394 1356 -1048
rect 860 -1395 1356 -1394
rect 732 -1414 1356 -1395
rect 1446 -1414 2127 -1048
rect 2208 -1213 2393 -893
rect 732 -1438 2127 -1414
rect 2209 -1402 2393 -1213
rect 732 -2094 891 -1438
rect 1623 -1579 1679 -1572
rect 1623 -1845 1679 -1639
rect 1043 -1901 1051 -1845
rect 1128 -1901 1728 -1845
rect 1805 -1901 1816 -1845
rect 2209 -2026 2217 -1402
rect 2387 -2026 2393 -1402
rect 732 -2113 2110 -2094
rect 732 -2118 2122 -2113
rect 732 -2255 746 -2118
rect 850 -2255 973 -2118
rect 1077 -2128 2122 -2118
rect 1077 -2252 1329 -2128
rect 1434 -2252 2122 -2128
rect 1077 -2255 2122 -2252
rect 732 -2267 2122 -2255
rect 733 -2357 2122 -2328
rect 733 -2494 1172 -2357
rect 1276 -2494 1558 -2357
rect 1662 -2494 1756 -2357
rect 1860 -2494 1984 -2357
rect 2088 -2358 2122 -2357
rect 2209 -2358 2393 -2026
rect 2088 -2494 2393 -2358
rect 733 -2542 2393 -2494
rect 529 -2679 849 -2670
rect 529 -2898 542 -2679
rect 840 -2898 849 -2679
rect 529 -2905 849 -2898
use sky130_fd_pr__pfet_g5v0d10v5_GTJ6Y6  sky130_fd_pr__pfet_g5v0d10v5_GTJ6Y6_0 paramcells
timestamp 1718242007
transform 1 0 1585 0 -1 232
box -387 -512 387 512
use sky130_fd_pr__pfet_g5v0d10v5_U6NWY6  sky130_fd_pr__pfet_g5v0d10v5_U6NWY6_0 paramcells
timestamp 1718242347
transform 1 0 1427 0 1 -1038
box -387 -762 387 762
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  sky130_fd_pr__pfet_g5v0d10v5_U62SY6_0 paramcells
timestamp 1718242097
transform 1 0 1932 0 1 -1038
box -308 -762 308 762
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  sky130_fd_pr__pfet_g5v0d10v5_U62SY6_1
timestamp 1718242097
transform 1 0 922 0 1 -1038
box -308 -762 308 762
use sky130_fd_pr__diode_pw2nd_11v0_QK8PWZ  XD1 paramcells
timestamp 1750254798
transform 1 0 1987 0 1 1055
box -217 -217 217 217
use sky130_fd_pr__nfet_g5v0d10v5_EJGQFX  XM1 paramcells
timestamp 1718240546
transform -1 0 1417 0 1 -2308
box -357 -458 357 458
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM3 paramcells
timestamp 1718240546
transform -1 0 907 0 1 -2308
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM5
timestamp 1718240546
transform 1 0 1927 0 1 -2308
box -278 -458 278 458
use sky130_fd_pr__pfet_g5v0d10v5_GTJ6Y6  XM7
timestamp 1718242007
transform 1 0 1001 0 -1 232
box -387 -512 387 512
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM8
timestamp 1718240546
transform 1 0 964 0 -1 1296
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM10
timestamp 1718240546
transform 1 0 1546 0 -1 1296
box -278 -458 278 458
<< labels >>
flabel metal1 326 -352 526 -152 0 FreeSans 256 0 0 0 vdd
port 5 nsew
flabel metal1 1705 773 1705 773 0 FreeSans 320 0 0 0 holdp
flabel metal1 1271 778 1271 778 0 FreeSans 320 0 0 0 holdb
flabel metal1 336 -2891 536 -2691 0 FreeSans 256 0 0 0 vss
port 2 nsew
flabel metal1 2326 -1396 2526 -1196 0 FreeSans 256 0 0 0 out
port 3 nsew
flabel metal1 333 -1397 533 -1197 0 FreeSans 256 0 0 0 in
port 4 nsew
flabel metal1 340 790 540 990 0 FreeSans 256 0 0 0 hold
port 1 nsew
<< end >>
