** sch_path: /home/tim/gits/chipalooza_projects_2/dependencies/sky130_ef_ip__samplehold/xschem/sky130_ef_ip__samplehold.sch
.subckt sky130_ef_ip__samplehold dvdd dvss hold vdd out in ena vss
*.PININFO vdd:I hold:I in:I vss:I out:O dvdd:I dvss:I ena:I
XC1 holdval vss sky130_fd_pr__cap_mim_m3_1 W=5 L=5 m=48
XC2 vss holdval sky130_fd_pr__cap_mim_m3_2 W=5 L=5 m=48
x1 hold3v vss holdval net1 vdd balanced_switch
x2 vdd out ena3v vss holdval dvss follower_amp
x3 vdd net1 ena3v vss in dvss follower_amp
x4 hold dvdd dvss dvss vdd vdd hold3v sky130_fd_sc_hvl__lsbuflv2hv_1
XXD1 dvss hold sky130_fd_pr__diode_pw2nd_05v5 area=3.6e11 perim=2.4e6
x5 ena dvdd dvss dvss vdd vdd ena3v sky130_fd_sc_hvl__lsbuflv2hv_1
XXD2 dvss ena sky130_fd_pr__diode_pw2nd_05v5 area=3.6e11 perim=2.4e6
.ends

* expanding   symbol:  balanced_switch.sym # of pins=5
** sym_path: /home/tim/gits/chipalooza_projects_2/dependencies/sky130_ef_ip__samplehold/xschem/balanced_switch.sym
** sch_path: /home/tim/gits/chipalooza_projects_2/dependencies/sky130_ef_ip__samplehold/xschem/balanced_switch.sch
.subckt balanced_switch hold vss out in vdd
*.PININFO in:I out:O vss:I vdd:I hold:I
XM1 in holdb out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
XM2 in holdp out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=2 m=1
XM3 out holdp out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM4 out holdb out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM5 in holdp in vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM6 in holdb in vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM7 holdb hold vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM8 holdb hold vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM9 holdp holdb vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 nf=1 m=1
XM10 holdp holdb vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XXD1 vss hold sky130_fd_pr__diode_pw2nd_11v0 area=2.025e11 perim=1.8e6
.ends


* expanding   symbol:  follower_amp.sym # of pins=6
** sym_path: /home/tim/gits/chipalooza_projects_2/dependencies/sky130_ef_ip__samplehold/xschem/follower_amp.sym
** sch_path: /home/tim/gits/chipalooza_projects_2/dependencies/sky130_ef_ip__samplehold/xschem/follower_amp.sch
.subckt follower_amp vdd out ena vss in vsub
*.PININFO in:I vdd:I vss:I out:O ena:I vsub:I
XM4 pdrv1 net1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM5 vdd net1 net1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM10 vss nbias nbias vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM20 out pdrv1 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=280 nf=280 m=1
XM22 out ndrv vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=4 m=1
XM24 pbias nbias vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM25 vdd pbias pbias vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM26 vcomp pbias vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM27 net2 out vcomp vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM28 vcomp in ndrv vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM29 ndrv net2 vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM30 vss net2 net2 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM1 net1 out vcomn1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM2 vcomn1 in pdrv1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM3 pdrv2 net3 vdd vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM6 vdd net3 net3 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM7 vcomn2 nbias vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM12 vdd pdrv2 out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=20 nf=20 m=1
XXD1 vss in sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
XM13 net4 ena nbias vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XXD2 vss ena sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
XM11 pdrv2 in vcomn2 vss sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 m=1
XM9 net3 out vcomn2 vss sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 m=1
XM8 vcomn1 nbias vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XR2 net4 vdd vss sky130_fd_pr__res_xhigh_po_0p35 L=140 mult=1 m=1
.ends

