magic
tech sky130A
magscale 1 2
timestamp 1740448282
<< locali >>
rect 813 10343 1130 10366
rect 813 10186 836 10343
rect 1105 10186 1130 10343
rect 813 10151 1130 10186
rect 938 9528 1068 10151
rect 557 9209 837 9231
rect 557 9120 575 9209
rect 818 9120 837 9209
rect 557 9097 837 9120
rect 2398 8510 2507 8539
rect 2398 8101 2414 8510
rect 2483 8101 2507 8510
rect 2398 8077 2507 8101
rect 2401 7685 2504 7713
rect 2401 7276 2418 7685
rect 2487 7276 2504 7685
rect 2401 7252 2504 7276
rect 557 6697 837 6721
rect 557 6608 576 6697
rect 819 6608 837 6697
rect 557 6587 837 6608
rect 975 5851 1105 6294
rect 814 5813 1131 5851
rect 814 5601 841 5813
rect 1098 5601 1131 5813
rect 814 5574 1131 5601
<< viali >>
rect 836 10186 1105 10343
rect 575 9120 818 9209
rect 2414 8101 2483 8510
rect 2418 7276 2487 7685
rect 576 6608 819 6697
rect 841 5601 1098 5813
<< metal1 >>
rect 134 11209 15840 11255
rect 134 10961 15354 11209
rect 134 10514 1726 10961
rect 2238 10538 15354 10961
rect 15799 10538 15840 11209
rect 2238 10514 15840 10538
rect 134 10494 15840 10514
rect 813 10343 3274 10367
rect 813 10186 836 10343
rect 1105 10260 3274 10343
rect 1105 10186 1130 10260
rect 813 10151 1130 10186
rect 2763 10024 3105 10046
rect 785 9713 831 10014
rect 241 9667 831 9713
rect 2763 9706 2783 10024
rect 3086 9706 3105 10024
rect 241 9255 287 9667
rect 338 9545 2459 9547
rect 338 9438 831 9545
rect 1122 9438 2459 9545
rect 52 9197 287 9255
rect 557 9209 837 9231
rect 557 9197 575 9209
rect 52 9128 575 9197
rect 52 9055 249 9128
rect 557 9120 575 9128
rect 818 9120 837 9209
rect 557 9097 837 9120
rect 2763 8848 3105 9706
rect 141 8834 688 8848
rect 2433 8834 3105 8848
rect 141 8824 3105 8834
rect 141 8564 167 8824
rect 663 8618 3105 8824
rect 663 8564 688 8618
rect 2433 8598 3105 8618
rect 141 8539 688 8564
rect 2398 8510 2507 8539
rect 2398 8101 2414 8510
rect 2483 8127 2507 8510
rect 2483 8101 2651 8127
rect 2398 8077 2651 8101
rect 2445 8076 2651 8077
rect 337 8001 2445 8010
rect 337 7796 831 8001
rect 1113 7796 2445 8001
rect 337 7794 2445 7796
rect 2401 7685 2550 7713
rect 148 7262 689 7292
rect 148 6997 171 7262
rect 662 7208 689 7262
rect 2401 7276 2418 7685
rect 2487 7276 2550 7685
rect 2401 7252 2550 7276
rect 662 6997 2448 7208
rect 148 6992 2448 6997
rect 148 6973 689 6992
rect 1263 6941 1581 6942
rect 1263 6867 1271 6941
rect 1571 6867 1581 6941
rect 1263 6855 1581 6867
rect 52 6686 252 6739
rect 557 6697 837 6721
rect 557 6686 576 6697
rect 52 6617 576 6686
rect 52 6539 287 6617
rect 557 6608 576 6617
rect 819 6608 837 6697
rect 557 6587 837 6608
rect 238 6140 287 6539
rect 341 6262 827 6393
rect 1123 6262 2447 6393
rect 341 6260 2447 6262
rect 1727 6151 2222 6193
rect 238 6091 855 6140
rect 806 5926 855 6091
rect 814 5851 855 5852
rect 814 5813 1131 5851
rect 814 5601 841 5813
rect 1098 5601 1131 5813
rect 1727 5823 1772 6151
rect 2178 5823 2222 6151
rect 1727 5645 2222 5823
rect 814 5574 1131 5601
rect 1725 5634 2222 5645
rect 1725 5367 2221 5634
rect 2501 5173 2550 7252
rect 2600 6556 2651 8076
rect 2600 6457 2654 6556
rect 2600 5153 2651 6457
rect 2763 5866 3105 8598
rect 2763 5833 15760 5866
rect 2763 5252 8148 5833
rect 8752 5286 11370 5833
rect 11984 5819 15760 5833
rect 11984 5286 14806 5819
rect 8752 5272 14806 5286
rect 15420 5272 15760 5819
rect 8752 5252 15760 5272
rect 2763 5224 15760 5252
rect 2193 3676 2906 3876
rect 3106 3676 3113 3876
rect 167 2559 623 2588
rect 167 1838 201 2559
rect 590 1838 623 2559
rect 167 1796 623 1838
rect 2172 1621 2504 1691
rect 2328 895 2681 914
rect 2328 709 2340 895
rect 2667 852 2681 895
rect 2667 738 3263 852
rect 2667 709 2681 738
rect 2328 679 2681 709
rect 2405 590 15829 630
rect 2405 585 14809 590
rect 2405 579 11370 585
rect 2405 557 8119 579
rect 127 535 8119 557
rect 127 171 159 535
rect 665 201 8119 535
rect 8706 207 11370 579
rect 11957 212 14809 585
rect 15396 212 15829 590
rect 11957 207 15829 212
rect 8706 201 15829 207
rect 665 171 15829 201
rect 127 153 15829 171
<< via1 >>
rect 1726 10514 2238 10961
rect 15354 10538 15799 11209
rect 836 10186 1105 10343
rect 2783 9706 3086 10024
rect 831 9423 1122 9545
rect 1271 8876 1573 8933
rect 167 8564 663 8824
rect 831 7796 1113 8001
rect 171 6997 662 7262
rect 1271 6867 1571 6941
rect 827 6262 1123 6394
rect 841 5601 1098 5813
rect 1772 5823 2178 6151
rect 8148 5252 8752 5833
rect 11370 5286 11984 5833
rect 14806 5272 15420 5819
rect 2906 3676 3106 3876
rect 201 1838 590 2559
rect 2340 709 2667 895
rect 159 171 665 535
rect 8119 201 8706 579
rect 11370 207 11957 585
rect 14809 212 15396 590
<< metal2 >>
rect 1702 10961 2256 10982
rect 1702 10514 1726 10961
rect 2238 10514 2256 10961
rect 1702 10494 2256 10514
rect 813 10343 1130 10366
rect 813 10186 836 10343
rect 1105 10186 1130 10343
rect 813 10151 1130 10186
rect 7578 10076 7778 11249
rect 15327 11209 15837 11245
rect 15327 10538 15354 11209
rect 15799 10538 15837 11209
rect 15327 10506 15837 10538
rect 143 10024 3111 10040
rect 143 9806 2783 10024
rect 143 9723 169 9806
rect 649 9723 2783 9806
rect 143 9706 2783 9723
rect 3086 9706 3111 10024
rect 143 9689 3111 9706
rect 813 9583 1136 9600
rect 813 9376 831 9583
rect 1122 9376 1136 9583
rect 813 9359 1136 9376
rect 1263 9011 1582 9021
rect 1263 8933 1272 9011
rect 1263 8876 1271 8933
rect 1574 8889 1582 9011
rect 1573 8876 1582 8889
rect 141 8824 688 8848
rect 141 8564 167 8824
rect 663 8564 688 8824
rect 141 8539 688 8564
rect 816 8029 1132 8042
rect 816 7796 831 8029
rect 1113 7796 1132 8029
rect 816 7771 1132 7796
rect 148 7262 689 7292
rect 148 6997 171 7262
rect 662 6997 689 7262
rect 148 6973 689 6997
rect 1263 6941 1582 6942
rect 1263 6746 1271 6941
rect 1571 6867 1582 6941
rect 1570 6746 1582 6867
rect 1263 6736 1582 6746
rect 2598 6461 2602 6506
rect 813 6430 1130 6442
rect 813 6394 828 6430
rect 1118 6394 1130 6430
rect 813 6262 827 6394
rect 1123 6262 1130 6394
rect 813 6234 828 6262
rect 1118 6234 1130 6262
rect 2654 6261 6128 6306
rect 813 6217 1130 6234
rect 1727 6152 2222 6193
rect 6421 6152 6939 6346
rect 1727 6151 6939 6152
rect 814 5813 1131 5851
rect 814 5601 841 5813
rect 1098 5601 1131 5813
rect 1727 5823 1772 6151
rect 2178 5823 6939 6151
rect 1727 5689 1775 5823
rect 2175 5689 6939 5823
rect 1727 5634 6939 5689
rect 814 5574 1131 5601
rect 1407 5467 2587 5596
rect 7660 5467 7860 6266
rect 1407 5456 7860 5467
rect 1407 5414 2839 5456
rect 1407 5001 1592 5414
rect 2369 5295 2839 5414
rect 3202 5295 7860 5456
rect 2369 5282 7860 5295
rect 8106 5892 8594 6322
rect 8106 5833 8791 5892
rect 8106 5252 8148 5833
rect 8752 5252 8791 5833
rect 11335 5884 11785 6352
rect 11335 5833 12020 5884
rect 15056 5871 15458 6337
rect 11335 5286 11370 5833
rect 11984 5286 12020 5833
rect 11335 5254 12020 5286
rect 14773 5819 15458 5871
rect 14773 5272 14806 5819
rect 15420 5272 15458 5819
rect 8106 5224 8791 5252
rect 14773 5239 15458 5272
rect 167 2559 623 2588
rect 167 1838 201 2559
rect 590 1838 623 2559
rect 2508 1885 2552 4984
rect 167 1796 623 1838
rect 2603 1004 2653 5134
rect 2906 4973 6390 5173
rect 2906 3876 3106 4973
rect 6190 4806 6390 4973
rect 2906 3667 3106 3676
rect 2603 954 6124 1004
rect 2328 895 2681 914
rect 2328 709 2340 895
rect 2667 709 2681 895
rect 2328 694 2681 709
rect 6422 654 6940 1065
rect 138 623 687 649
rect 138 171 159 623
rect 665 171 687 623
rect 2187 549 6940 654
rect 138 149 687 171
rect 1684 508 6940 549
rect 1684 165 1727 508
rect 2235 165 6940 508
rect 1684 136 6940 165
rect 7661 119 7861 1001
rect 8070 654 8557 1067
rect 8070 579 8755 654
rect 11476 646 11863 1109
rect 15057 663 15441 1070
rect 8070 201 8119 579
rect 8706 201 8755 579
rect 8070 154 8755 201
rect 11316 585 12001 646
rect 11316 207 11370 585
rect 11957 207 12001 585
rect 11316 157 12001 207
rect 14756 590 15441 663
rect 14756 212 14809 590
rect 15396 212 15441 590
rect 14756 157 15441 212
<< via2 >>
rect 1726 10514 2238 10961
rect 836 10186 1105 10343
rect 15354 10538 15799 11209
rect 169 9723 649 9806
rect 831 9545 1122 9583
rect 831 9423 1122 9545
rect 831 9376 1122 9423
rect 1272 8933 1574 9011
rect 1272 8889 1573 8933
rect 1573 8889 1574 8933
rect 167 8564 663 8824
rect 831 8001 1113 8029
rect 831 7796 1113 8001
rect 171 6997 662 7262
rect 1271 6867 1570 6930
rect 1271 6746 1570 6867
rect 828 6394 1118 6430
rect 828 6262 1118 6394
rect 828 6234 1118 6262
rect 841 5601 1098 5813
rect 1775 5823 2175 6140
rect 1775 5689 2175 5823
rect 2839 5295 3202 5456
rect 201 1838 590 2559
rect 2340 709 2667 895
rect 159 535 665 623
rect 159 171 665 535
rect 1727 165 2235 508
<< metal3 >>
rect 133 11046 694 11255
rect 813 11046 1133 11254
rect 1263 11250 1582 11253
rect 1263 11048 1583 11250
rect 138 9806 692 11046
rect 138 9723 169 9806
rect 649 9723 692 9806
rect 138 8824 692 9723
rect 138 8564 167 8824
rect 663 8564 692 8824
rect 138 7262 692 8564
rect 138 6997 171 7262
rect 662 6997 692 7262
rect 138 2559 692 6997
rect 138 1838 201 2559
rect 590 1838 692 2559
rect 138 1289 692 1838
rect 813 10343 1132 11046
rect 813 10186 836 10343
rect 1105 10186 1132 10343
rect 813 9583 1132 10186
rect 813 9376 831 9583
rect 1122 9376 1132 9583
rect 813 8029 1132 9376
rect 813 7796 831 8029
rect 1113 7796 1132 8029
rect 813 6430 1132 7796
rect 813 6234 828 6430
rect 1118 6234 1132 6430
rect 813 5813 1132 6234
rect 813 5601 841 5813
rect 1098 5601 1132 5813
rect 138 623 687 1289
rect 138 171 159 623
rect 665 171 687 623
rect 138 0 687 171
rect 813 943 1132 5601
rect 813 674 840 943
rect 1101 674 1132 943
rect 813 0 1132 674
rect 1263 9011 1582 11048
rect 1263 8889 1272 9011
rect 1574 8889 1582 9011
rect 1263 6930 1582 8889
rect 1263 6746 1271 6930
rect 1570 6746 1582 6930
rect 1263 0 1582 6746
rect 1702 10961 2256 11253
rect 1702 10514 1726 10961
rect 2238 10514 2256 10961
rect 1702 6215 2256 10514
rect 15327 11209 15837 11245
rect 15327 10538 15354 11209
rect 15799 10538 15837 11209
rect 15327 10506 15837 10538
rect 1692 6140 2256 6215
rect 1692 5689 1775 6140
rect 2175 5689 2256 6140
rect 1692 5621 2256 5689
rect 1702 508 2256 5621
rect 2821 5475 3216 5494
rect 2821 5242 2838 5475
rect 3196 5456 3216 5475
rect 3202 5295 3216 5456
rect 3196 5242 3216 5295
rect 2821 5225 3216 5242
rect 2328 895 2681 914
rect 2328 709 2340 895
rect 2667 709 2681 895
rect 2328 679 2681 709
rect 1702 165 1727 508
rect 2235 165 2256 508
rect 1702 0 2256 165
<< via3 >>
rect 840 674 1101 943
rect 15354 10538 15799 11209
rect 2838 5456 3196 5475
rect 2838 5295 2839 5456
rect 2839 5295 3196 5456
rect 2838 5242 3196 5295
rect 2340 709 2667 895
<< metal4 >>
rect 13833 11209 15845 11245
rect 13833 10538 15354 11209
rect 15799 10538 15845 11209
rect 13833 10506 15845 10538
rect 2813 5546 3228 5576
rect 2813 5213 2838 5546
rect 2814 4653 2838 5213
rect 3196 4653 3228 5546
rect 2814 4624 3228 4653
rect 813 943 2683 970
rect 813 674 840 943
rect 1101 895 2683 943
rect 1101 709 2340 895
rect 2667 709 2683 895
rect 1101 674 2683 709
rect 813 651 2683 674
<< via4 >>
rect 2838 5475 3196 5546
rect 2838 5242 3196 5475
rect 2838 4653 3196 5242
<< metal5 >>
rect 2813 5546 3228 5576
rect 2813 5213 2838 5546
rect 2814 4653 2838 5213
rect 3196 4653 3228 5546
rect 2814 4624 3228 4653
use amp_via_4cut  amp_via_4cut_0
timestamp 1718240546
transform 0 1 10525 -1 0 21136
box 15948 -7932 16222 -7868
use amp_via_4cut  amp_via_4cut_1
timestamp 1718240546
transform 0 1 10528 -1 0 22473
box 15948 -7932 16222 -7868
use amp_via_4cut  amp_via_4cut_2
timestamp 1718240546
transform 0 1 10425 -1 0 21136
box 15948 -7932 16222 -7868
use amp_via_4cut  amp_via_4cut_3
timestamp 1718240546
transform 0 1 10430 -1 0 17839
box 15948 -7932 16222 -7868
use hold_cap_array  hold_cap_array_0
timestamp 1718240546
transform 0 1 29374 -1 0 13175
box 1925 -26553 13175 -15183
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_0 paramcells
timestamp 1718240546
transform 1 0 849 0 1 5980
box -198 -198 198 198
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_1
timestamp 1718240546
transform 1 0 814 0 1 10008
box -198 -198 198 198
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1738263620
transform 1 0 338 0 -1 9537
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_1
timestamp 1738263620
transform 1 0 338 0 1 6281
box -66 -43 2178 1671
use balanced_switch  x1
timestamp 1719257891
transform -1 0 2543 0 -1 2480
box 301 -3111 2543 2130
use follower_amp  x2
timestamp 1740434940
transform 0 1 4681 1 0 743
box 0 -1436 4377 11129
use follower_amp  x3
timestamp 1740434940
transform 0 1 4680 1 0 5991
box 0 -1436 4377 11129
<< labels >>
flabel metal3 1703 11046 2255 11253 0 FreeSans 1600 90 0 0 vss
port 5 nsew
flabel metal3 1263 11048 1583 11250 0 FreeSans 1600 90 0 0 dvdd
port 6 nsew
flabel metal3 813 11046 1133 11254 0 FreeSans 1600 90 0 0 dvss
port 7 nsew
flabel metal3 133 11046 694 11255 0 FreeSans 1600 90 0 0 vdd
port 2 nsew
flabel metal1 52 9055 249 9255 0 FreeSans 320 0 0 0 ena
port 8 nsew
flabel metal1 52 6539 252 6739 0 FreeSans 256 0 0 0 hold
port 3 nsew
flabel metal2 7661 119 7861 319 0 FreeSans 256 0 0 0 in
port 4 nsew
flabel metal2 7578 11049 7778 11249 0 FreeSans 256 270 0 0 out
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 15845 11255
<< end >>
