magic
tech sky130A
magscale 1 2
timestamp 1750254930
<< locali >>
rect 813 10343 1130 10366
rect 813 10186 836 10343
rect 1105 10186 1130 10343
rect 813 10151 1130 10186
rect 938 9528 1068 10151
rect 557 9209 837 9231
rect 557 9120 575 9209
rect 818 9120 837 9209
rect 557 9097 837 9120
rect 2398 8510 2507 8539
rect 2398 8101 2414 8510
rect 2483 8101 2507 8510
rect 2398 8077 2507 8101
rect 2401 7685 2504 7713
rect 2401 7276 2418 7685
rect 2487 7276 2504 7685
rect 2401 7252 2504 7276
rect 557 6697 837 6721
rect 557 6608 576 6697
rect 819 6608 837 6697
rect 557 6587 837 6608
rect 975 5851 1105 6294
rect 814 5813 1131 5851
rect 814 5601 841 5813
rect 1098 5601 1131 5813
rect 814 5574 1131 5601
<< viali >>
rect 836 10186 1105 10343
rect 575 9120 818 9209
rect 2414 8101 2483 8510
rect 2418 7276 2487 7685
rect 576 6608 819 6697
rect 841 5601 1098 5813
<< metal1 >>
rect 134 11209 15901 11255
rect 134 10961 15415 11209
rect 134 10514 1726 10961
rect 2238 10538 15415 10961
rect 15860 10538 15901 11209
rect 2238 10537 15901 10538
rect 2238 10514 3080 10537
rect 134 10494 3080 10514
rect 813 10343 3300 10367
rect 813 10186 836 10343
rect 1105 10260 3300 10343
rect 1105 10186 1130 10260
rect 813 10151 1130 10186
rect 2824 10024 3166 10046
rect 785 9713 831 10014
rect 241 9667 831 9713
rect 2824 9706 2844 10024
rect 3147 9706 3166 10024
rect 241 9255 287 9667
rect 338 9545 2459 9547
rect 338 9438 831 9545
rect 1122 9438 2459 9545
rect 52 9197 287 9255
rect 557 9209 837 9231
rect 557 9197 575 9209
rect 52 9128 575 9197
rect 52 9055 249 9128
rect 557 9120 575 9128
rect 818 9120 837 9209
rect 557 9097 837 9120
rect 2824 8848 3166 9706
rect 141 8834 688 8848
rect 2433 8834 3166 8848
rect 141 8824 3166 8834
rect 141 8564 167 8824
rect 663 8618 3166 8824
rect 663 8564 688 8618
rect 2433 8598 3166 8618
rect 141 8539 688 8564
rect 2398 8510 2507 8539
rect 2398 8101 2414 8510
rect 2483 8127 2507 8510
rect 2483 8101 2651 8127
rect 2398 8077 2651 8101
rect 2445 8076 2651 8077
rect 337 8001 2445 8010
rect 337 7796 831 8001
rect 1113 7796 2445 8001
rect 337 7794 2445 7796
rect 2401 7685 2550 7713
rect 148 7262 689 7292
rect 148 6997 171 7262
rect 662 7208 689 7262
rect 2401 7276 2418 7685
rect 2487 7276 2550 7685
rect 2401 7252 2550 7276
rect 662 6997 2448 7208
rect 148 6992 2448 6997
rect 148 6973 689 6992
rect 1263 6941 1581 6942
rect 1263 6867 1271 6941
rect 1571 6867 1581 6941
rect 1263 6855 1581 6867
rect 52 6686 252 6739
rect 557 6697 837 6721
rect 557 6686 576 6697
rect 52 6617 576 6686
rect 52 6539 287 6617
rect 557 6608 576 6617
rect 819 6608 837 6697
rect 557 6587 837 6608
rect 238 6140 287 6539
rect 341 6262 827 6393
rect 1123 6262 2447 6393
rect 341 6260 2447 6262
rect 1727 6151 2222 6193
rect 238 6091 855 6140
rect 806 5926 855 6091
rect 814 5851 855 5852
rect 814 5813 1131 5851
rect 814 5601 841 5813
rect 1098 5601 1131 5813
rect 1727 5823 1772 6151
rect 2178 5823 2222 6151
rect 1727 5645 2222 5823
rect 814 5574 1131 5601
rect 1725 5634 2222 5645
rect 1725 5367 2221 5634
rect 2501 5173 2550 7252
rect 2600 6556 2651 8076
rect 2600 6457 2654 6556
rect 2600 5153 2651 6457
rect 2824 5866 3166 8598
rect 2824 5833 15821 5866
rect 2824 5271 8209 5833
rect 8813 5286 11431 5833
rect 12045 5819 15821 5833
rect 12045 5286 14867 5819
rect 8813 5272 14867 5286
rect 15481 5272 15821 5819
rect 8813 5271 15821 5272
rect 2193 3676 2962 3876
rect 3162 3676 3169 3876
rect 167 2559 623 2588
rect 167 1838 201 2559
rect 590 1838 623 2559
rect 167 1796 623 1838
rect 2172 1621 2504 1691
rect 2328 895 2681 914
rect 2328 709 2340 895
rect 2667 852 2681 895
rect 2667 738 3324 852
rect 2667 709 2681 738
rect 2328 679 2681 709
rect 2405 590 15890 630
rect 2405 585 14870 590
rect 2405 579 11431 585
rect 2405 557 8180 579
rect 127 535 8180 557
rect 127 171 159 535
rect 665 201 8180 535
rect 8767 207 11431 579
rect 12018 212 14870 585
rect 15457 212 15890 590
rect 12018 207 15890 212
rect 8767 201 15890 207
rect 665 171 15890 201
rect 127 153 15890 171
<< via1 >>
rect 1726 10514 2238 10961
rect 15415 10538 15860 11209
rect 836 10186 1105 10343
rect 2844 9706 3147 10024
rect 831 9423 1122 9545
rect 1271 8876 1573 8933
rect 167 8564 663 8824
rect 831 7796 1113 8001
rect 171 6997 662 7262
rect 1271 6867 1571 6941
rect 827 6262 1123 6394
rect 841 5601 1098 5813
rect 1772 5823 2178 6151
rect 8209 5271 8813 5833
rect 11431 5286 12045 5833
rect 14867 5272 15481 5819
rect 2962 3676 3162 3876
rect 201 1838 590 2559
rect 2340 709 2667 895
rect 159 171 665 535
rect 8180 201 8767 579
rect 11431 207 12018 585
rect 14870 212 15457 590
<< metal2 >>
rect 1702 10961 2256 10982
rect 1702 10514 1726 10961
rect 2238 10514 2256 10961
rect 1702 10494 2256 10514
rect 813 10343 1130 10366
rect 813 10186 836 10343
rect 1105 10186 1130 10343
rect 813 10151 1130 10186
rect 7639 10076 7839 11249
rect 15388 11209 15898 11245
rect 15388 10538 15415 11209
rect 15860 10538 15898 11209
rect 15388 10506 15898 10538
rect 143 10024 3172 10040
rect 143 9806 2844 10024
rect 143 9723 169 9806
rect 649 9723 2844 9806
rect 143 9706 2844 9723
rect 3147 9706 3172 10024
rect 143 9689 3172 9706
rect 813 9583 1136 9600
rect 813 9376 831 9583
rect 1122 9376 1136 9583
rect 813 9359 1136 9376
rect 1263 9011 1582 9021
rect 1263 8933 1272 9011
rect 1263 8876 1271 8933
rect 1574 8889 1582 9011
rect 1573 8876 1582 8889
rect 141 8824 688 8848
rect 141 8564 167 8824
rect 663 8564 688 8824
rect 141 8539 688 8564
rect 816 8029 1132 8042
rect 816 7796 831 8029
rect 1113 7796 1132 8029
rect 816 7771 1132 7796
rect 148 7262 689 7292
rect 148 6997 171 7262
rect 662 6997 689 7262
rect 148 6973 689 6997
rect 1263 6941 1582 6942
rect 1263 6746 1271 6941
rect 1571 6867 1582 6941
rect 1570 6746 1582 6867
rect 1263 6736 1582 6746
rect 2598 6461 2602 6506
rect 813 6430 1130 6442
rect 813 6394 828 6430
rect 1118 6394 1130 6430
rect 813 6262 827 6394
rect 1123 6262 1130 6394
rect 813 6234 828 6262
rect 1118 6234 1130 6262
rect 2654 6261 6189 6306
rect 813 6217 1130 6234
rect 1727 6152 2222 6193
rect 6482 6152 7000 6346
rect 1727 6151 7000 6152
rect 814 5813 1131 5851
rect 814 5601 841 5813
rect 1098 5601 1131 5813
rect 1727 5823 1772 6151
rect 2178 5823 7000 6151
rect 1727 5689 1775 5823
rect 2175 5689 7000 5823
rect 1727 5634 7000 5689
rect 814 5574 1131 5601
rect 1407 5547 2587 5596
rect 7721 5547 7921 6269
rect 1407 5536 7921 5547
rect 1407 5414 2900 5536
rect 1407 5001 1592 5414
rect 2369 5375 2900 5414
rect 3263 5375 7921 5536
rect 2369 5362 7921 5375
rect 8167 5892 8655 6322
rect 8167 5833 8852 5892
rect 8167 5271 8209 5833
rect 8813 5271 8852 5833
rect 167 2559 623 2588
rect 167 1838 201 2559
rect 590 1838 623 2559
rect 2508 1885 2552 4984
rect 167 1796 623 1838
rect 2603 1004 2653 5134
rect 2962 5072 6484 5268
rect 8167 5224 8852 5271
rect 11396 5884 11846 6352
rect 11396 5833 12081 5884
rect 15117 5871 15519 6337
rect 11396 5286 11431 5833
rect 12045 5286 12081 5833
rect 11396 5254 12081 5286
rect 14834 5819 15519 5871
rect 14834 5272 14867 5819
rect 15481 5272 15519 5819
rect 14834 5239 15519 5272
rect 2962 3876 3162 5072
rect 6252 4988 6484 5072
rect 2962 3667 3162 3676
rect 2603 954 6185 1004
rect 2328 895 2681 914
rect 2328 709 2340 895
rect 2667 709 2681 895
rect 2328 694 2681 709
rect 6483 654 7001 1065
rect 138 623 687 649
rect 138 171 159 623
rect 665 171 687 623
rect 2187 549 7001 654
rect 138 149 687 171
rect 1684 508 7001 549
rect 1684 165 1727 508
rect 2235 165 7001 508
rect 1684 136 7001 165
rect 7722 119 7922 1001
rect 8131 654 8618 1067
rect 8131 579 8816 654
rect 11537 646 11924 1109
rect 15118 663 15502 1070
rect 8131 201 8180 579
rect 8767 201 8816 579
rect 8131 154 8816 201
rect 11377 585 12062 646
rect 11377 207 11431 585
rect 12018 207 12062 585
rect 11377 157 12062 207
rect 14817 590 15502 663
rect 14817 212 14870 590
rect 15457 212 15502 590
rect 14817 157 15502 212
<< via2 >>
rect 1726 10514 2238 10961
rect 836 10186 1105 10343
rect 15415 10538 15860 11209
rect 169 9723 649 9806
rect 831 9545 1122 9583
rect 831 9423 1122 9545
rect 831 9376 1122 9423
rect 1272 8933 1574 9011
rect 1272 8889 1573 8933
rect 1573 8889 1574 8933
rect 167 8564 663 8824
rect 831 8001 1113 8029
rect 831 7796 1113 8001
rect 171 6997 662 7262
rect 1271 6867 1570 6930
rect 1271 6746 1570 6867
rect 828 6394 1118 6430
rect 828 6262 1118 6394
rect 828 6234 1118 6262
rect 841 5601 1098 5813
rect 1775 5823 2175 6140
rect 1775 5689 2175 5823
rect 2900 5375 3263 5536
rect 201 1838 590 2559
rect 2340 709 2667 895
rect 159 535 665 623
rect 159 171 665 535
rect 1727 165 2235 508
<< metal3 >>
rect 133 11046 694 11255
rect 813 11046 1133 11254
rect 1263 11250 1582 11253
rect 1263 11048 1583 11250
rect 138 9806 692 11046
rect 138 9723 169 9806
rect 649 9723 692 9806
rect 138 8824 692 9723
rect 138 8564 167 8824
rect 663 8564 692 8824
rect 138 7262 692 8564
rect 138 6997 171 7262
rect 662 6997 692 7262
rect 138 2559 692 6997
rect 138 1838 201 2559
rect 590 1838 692 2559
rect 138 1289 692 1838
rect 813 10343 1132 11046
rect 813 10186 836 10343
rect 1105 10186 1132 10343
rect 813 9583 1132 10186
rect 813 9376 831 9583
rect 1122 9376 1132 9583
rect 813 8029 1132 9376
rect 813 7796 831 8029
rect 1113 7796 1132 8029
rect 813 6430 1132 7796
rect 813 6234 828 6430
rect 1118 6234 1132 6430
rect 813 5813 1132 6234
rect 813 5601 841 5813
rect 1098 5601 1132 5813
rect 138 623 687 1289
rect 138 171 159 623
rect 665 171 687 623
rect 138 0 687 171
rect 813 943 1132 5601
rect 813 674 840 943
rect 1101 674 1132 943
rect 813 0 1132 674
rect 1263 9011 1582 11048
rect 1263 8889 1272 9011
rect 1574 8889 1582 9011
rect 1263 6930 1582 8889
rect 1263 6746 1271 6930
rect 1570 6746 1582 6930
rect 1263 0 1582 6746
rect 1702 10961 2256 11253
rect 1702 10514 1726 10961
rect 2238 10514 2256 10961
rect 1702 6215 2256 10514
rect 15388 11209 15898 11245
rect 15388 10538 15415 11209
rect 15860 10538 15898 11209
rect 15388 10506 15898 10538
rect 1692 6140 2256 6215
rect 1692 5689 1775 6140
rect 2175 5689 2256 6140
rect 1692 5621 2256 5689
rect 1702 508 2256 5621
rect 2882 5555 3277 5574
rect 2882 5242 2899 5555
rect 3257 5536 3277 5555
rect 3263 5375 3277 5536
rect 3257 5242 3277 5375
rect 2882 5225 3277 5242
rect 2328 895 2681 914
rect 2328 709 2340 895
rect 2667 709 2681 895
rect 2328 679 2681 709
rect 1702 165 1727 508
rect 2235 165 2256 508
rect 1702 0 2256 165
<< via3 >>
rect 840 674 1101 943
rect 15415 10538 15860 11209
rect 2899 5536 3257 5555
rect 2899 5375 2900 5536
rect 2900 5375 3257 5536
rect 2899 5242 3257 5375
rect 2340 709 2667 895
<< metal4 >>
rect 13894 11209 15906 11245
rect 13894 10538 15415 11209
rect 15860 10538 15906 11209
rect 13894 10506 15906 10538
rect 2874 5555 3289 5576
rect 2874 5213 2899 5555
rect 2875 4653 2899 5213
rect 3257 4653 3289 5555
rect 2875 4624 3289 4653
rect 813 943 2683 970
rect 813 674 840 943
rect 1101 895 2683 943
rect 1101 709 2340 895
rect 2667 709 2683 895
rect 1101 674 2683 709
rect 813 651 2683 674
<< via4 >>
rect 2899 5242 3257 5546
rect 2899 4653 3257 5242
<< metal5 >>
rect 2874 5546 3289 5576
rect 2874 5213 2899 5546
rect 2875 4653 2899 5213
rect 3257 4653 3289 5546
rect 2875 4624 3289 4653
use amp_via_4cut  amp_via_4cut_0
timestamp 1718240546
transform 0 1 10525 -1 0 21136
box 15948 -7932 16222 -7868
use amp_via_4cut  amp_via_4cut_1
timestamp 1718240546
transform 0 1 10528 -1 0 22473
box 15948 -7932 16222 -7868
use amp_via_4cut  amp_via_4cut_2
timestamp 1718240546
transform 0 1 10425 -1 0 21136
box 15948 -7932 16222 -7868
use amp_via_4cut  amp_via_4cut_3
timestamp 1718240546
transform 0 1 10430 -1 0 17839
box 15948 -7932 16222 -7868
use hold_cap_array  hold_cap_array_0
timestamp 1718240546
transform 0 1 29435 -1 0 13175
box 1925 -26553 13175 -15183
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_0 paramcells
timestamp 1718240546
transform 1 0 849 0 1 5980
box -198 -198 198 198
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_1
timestamp 1718240546
transform 1 0 814 0 1 10008
box -198 -198 198 198
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1750210935
transform 1 0 338 0 -1 9537
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_1
timestamp 1750210935
transform 1 0 338 0 1 6281
box -66 -43 2178 1671
use balanced_switch  x1
timestamp 1750254930
transform -1 0 2543 0 -1 2480
box 264 -3133 2570 2130
use follower_amp  x2
timestamp 1747667787
transform 0 1 4742 1 0 743
box 0 -1542 4469 11129
use follower_amp  x3
timestamp 1747667787
transform 0 1 4741 1 0 6011
box 0 -1542 4469 11129
<< labels >>
flabel metal3 1703 11046 2255 11253 0 FreeSans 1600 90 0 0 vss
port 5 nsew
flabel metal3 1263 11048 1583 11250 0 FreeSans 1600 90 0 0 dvdd
port 6 nsew
flabel metal3 813 11046 1133 11254 0 FreeSans 1600 90 0 0 dvss
port 7 nsew
flabel metal3 133 11046 694 11255 0 FreeSans 1600 90 0 0 vdd
port 2 nsew
flabel metal1 52 9055 249 9255 0 FreeSans 320 0 0 0 ena
port 8 nsew
flabel metal1 52 6539 252 6739 0 FreeSans 256 0 0 0 hold
port 3 nsew
flabel metal2 7722 119 7922 319 0 FreeSans 256 0 0 0 in
port 4 nsew
flabel metal2 7639 11049 7839 11249 0 FreeSans 256 270 0 0 out
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 15845 11255
<< end >>
